`timescale 1ns / 1ps
module counter(
    input       clk,
    input       areset,
    input       count_down_start,
    output reg [3:0] out_count_up,
    output reg [3:0] out_count_down
); 

    
//TODO


endmodule