`timescale 1ns / 1ps
module shift(
    input clk,      
    input [3:0] d,  
    input load,  
    output reg [3:0] q 
);

//TODO

endmodule