`timescale 1ns / 1ps
module flipflop (
    input clk,      
    input reset,   
    input d,       
    output reg q  
);

//TODO

endmodule