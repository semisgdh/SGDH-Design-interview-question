`timescale 1ns / 1ps
module fsm(
    input            clk,
    input            areset,
    input            in,
    output           out_fsm
); 

//TODO


endmodule