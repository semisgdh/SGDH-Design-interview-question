`timescale 1ns / 1ps
module basic_gate
(
    input in_a,
    input in_b,
    output not_gate_out,
    output and_gate_out,
    output nand_gate_out,
    output or_gate_out,
    output nor_gate_out,
    output xor_gate_out,
    output xnor_gate_out
);


//TODO


endmodule
