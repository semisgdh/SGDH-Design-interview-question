`timescale 1ns / 1ps
module module_top
(
input [1:0]     in_add_a,
input [1:0]     in_add_b,
input [1:0]     in_add_c,
input [1:0]     in_add_d,
input           in_add_sub_sel,
output [7:0]    final_cal_out

);

//TODO

endmodule
