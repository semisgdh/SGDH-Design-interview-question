`timescale 1ns / 1ps
module adder_position
(
input [1:0]     aklfjlskftnmnsfljksartnlkjhvlkjawlertkjdslgviuwelaktlsdhg,
input [1:0]     zkdjrhwekjtbmqiwuerbjcvmnxcvbksfjghoisogawtuhusguiuysadoi,
output [2:0]    klfgklrtlisrtgklbjkjkjilsdfljhsrgjkkjkjsdrtkukuhkukuhdrgk

);

assign klfgklrtlisrtgklbjkjkjilsdfljhsrgjkkjkjsdrtkukuhkukuhdrgk = aklfjlskftnmnsfljksartnlkjhvlkjawlertkjdslgviuwelaktlsdhg + zkdjrhwekjtbmqiwuerbjcvmnxcvbksfjghoisogawtuhusguiuysadoi;

endmodule
