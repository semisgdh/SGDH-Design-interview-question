`timescale 1ns / 1ps
module kmap
(
   input A,
   input B,
   input C,
   input D,
   output F_0,
   output F_1,
   output F_2
);

//#1 =====================================
//A B	C D  F_0 
//0 0	0 0   0
//0 0	0 1   1
//0 0	1 0   1
//0 0	1 1   0
//0 1	0 0   1
//0 1	0 1   0
//0 1	1 0   0
//0 1	1 1   1
//1 0	0 0   1
//1 0	0 1   0
//1 0	1 0   0
//1 0	1 1   1
//1 1	0 0   0
//1 1	0 1   1
//1 1	1 0   1
//1 1	1 1   0

//       CD
//    | 00 | 01 | 11 | 10 |
//   ----------------------
// AB |    |    |    |    |
// 00 |  0 |  1 |  0 |  1 |
// 01 |  1 |  0 |  1 |  0 |
// 11 |  0 |  1 |  0 |  1 |
// 10 |  1 |  0 |  1 |  0 |

// F = A'B'C'D + A'B'CD' + A'BC'D' + A'BCD + ABC'D + ABCD' + AB'C'D' + AB'CD

assign F_0 = (~A & ~B & ~C &  D) | 
             (~A & ~B &  C & ~D) |
             (~A &  B & ~C & ~D) |
             (~A &  B &  C &  D) |
             ( A &  B & ~C &  D) |
             ( A &  B &  C & ~D) |
             ( A & ~B & ~C & ~D) |
             ( A & ~B &  C &  D) ;
// #2 ==================================
// A	B	C	D	F_1
// 0	0	0	0	0
// 0	0	0	1	0
// 0	0	1	0	0
// 0	0	1	1	0
// 0	1	0	0	0
// 0	1	0	1	1
// 0	1	1	0	1
// 0	1	1	1	1
// 1	0	0	0	1
// 1	0	0	1	0
// 1	0	1	0	1
// 1	0	1	1	1
// 1	1	0	0	0
// 1	1	0	1	1
// 1	1	1	0	1
// 1	1	1	1	1
//       CD
//    | 00 | 01 | 11 | 10 |
//   ----------------------
// AB |    |    |    |    |
// 00 |  0 |  0 |  0 |  0 |
// 01 |  0 |  1 |  1 |  1 |
// 11 |  0 |  1 |  1 |  1 |
// 10 |  1 |  0 |  1 |  1 |
// F_1 = BD + BC + AC + AB'D'

assign F_1 = (B & D) | (B & C) | (A & C) | (A & ~B & ~D);

//#3=========================================
// A	B	C	D	F_2 돈케어 (X)
// 0	0	0	0	0	0
// 0	0	0	1	X	1
// 0	0	1	0	1	0
// 0	0	1	1	1	0
// 0	1	0	0	0	0
// 0	1	0	1	X	1
// 0	1	1	0	1	0
// 0	1	1	1	1	0
// 1	0	0	0	1	0
// 1	0	0	1	X	1
// 1	0	1	0	0	0
// 1	0	1	1	0	0
// 1	1	0	0	1	0
// 1	1	0	1	X	1
// 1	1	1	0	1	0
// 1	1	1	1	1	0
//        CD
//     | 00 | 01 | 11 | 10 |
//    ----------------------
//  AB |    |    |    |    |
//  00 |  0 |  X |  1 |  1 |
//  01 |  0 |  X |  1 |  1 |
//  11 |  1 |  X |  1 |  1 |
//  10 |  1 |  X |  0 |  0 |
// 
// F_2 = BC + A'C + AC'


assign F_2 = (B & C) | (~A & C) | (A & ~C);

endmodule
