`timescale 1ns / 1ps
module condition(
    input [1:0] sel,
    output reg [1:0] normal_if,   
    output reg [1:0] normal_case,   
    output     [1:0] normal_ternary,   
    output reg [1:0] latch_if,   
    output reg [1:0] latch_case   
); 

//TODO

endmodule